`include "TileAccumUnit/ReadPipeline/RemapCache/RemapCache.sv"
