`include "ParallelBlockLooper.sv"
