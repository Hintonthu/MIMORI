`include "TileAccumUnit/WritePipeline/WritePipeline.sv"
