`include "TileAccumUnit/AluPipeline/SimdDriver.sv"
