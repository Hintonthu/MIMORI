`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooper.sv"
