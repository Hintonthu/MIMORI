`include "TileAccumUnit/CoreAccumLooper.sv"
