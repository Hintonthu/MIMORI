`include "define.sv"
`include "common/ND.sv"
`include "common/BitOperation.sv"
`include "common/Controllers.sv"
`include "common/Registers.sv"
`include "common/OffsetStage.sv"
`include "TileAccumUnit/common/BofsExpand.sv"
`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooperIndexStage.sv"
`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooperStencilStage.sv"
`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooperMemofsStage.sv"
`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooperVectorStage.sv"
`include "TileAccumUnit/common/AccumWarpLooper.sv"
