`include "define.sv"
`include "TileAccumUnit/ReadPipeline/SramWriteCollector.sv"
