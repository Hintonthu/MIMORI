`include "TileAccumUnit/AccumBlockLooper.sv"
