`include "define.sv"
`include "TileAccumUnit/ReadPipeline/Allocator.sv"
