`include "TileAccumUnit/ReadPipeline/ReadPipeline.sv"
