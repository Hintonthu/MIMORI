`include "Top_mc.sv"
