`include "saed32sram.v"
`include "saed32nm.v"
`include "define.sv"
`include "TopGateWrap.sv"
`include "Top_syn.v"
