`include "common/SFifo.sv"
