`include "TileAccumUnit/ReadPipeline/SramWriteCollector.sv"
