`include "TileAccumUnit/TileAccumUnit.sv"
