`include "ParallelBlockLooper_sd.sv"
