`include "TileAccumUnit/DmaPipeline/DmaPipeline.sv"
