`include "define.sv"
`include "common/SRAM.sv"
`include "common/Controllers.sv"
`include "TileAccumUnit/ReadPipeline/RemapCache/BankSramReadIf.sv"
`include "TileAccumUnit/ReadPipeline/RemapCache/BankSramWriteButterflyIf.sv"
`include "TileAccumUnit/ReadPipeline/RemapCache/RemapCache.sv"
