`include "Top_sd.sv"
