`include "define.sv"
`include "common/ND.sv"
`include "common/BitOperation.sv"
`include "common/Controllers.sv"
`include "common/Registers.sv"
`include "common/OffsetStage.sv"
`include "common/SRAM.sv"
`include "common/IndexStage.sv"
`include "common/MemofsStage.sv"
`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooperCollector.sv"
`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooperIndexStage.sv"
`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooperStencilStage.sv"
`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooperMemofsStage.sv"
`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooperVectorStage.sv"
`include "TileAccumUnit/common/AccumWarpLooper.sv"
`include "TileAccumUnit/common/AccumBlockLooper.sv"
`include "TileAccumUnit/common/OrCrossBar.sv"
`include "TileAccumUnit/ReadPipeline/ChunkAddrLooper/ChunkRow.sv"
`include "TileAccumUnit/ReadPipeline/ChunkAddrLooper/ChunkRowStart.sv"
`include "TileAccumUnit/ReadPipeline/ChunkAddrLooper.sv"
`include "TileAccumUnit/ReadPipeline/RemapCache/BankSramReadIf.sv"
`include "TileAccumUnit/ReadPipeline/RemapCache/BankSramWriteButterflyIf.sv"
`include "TileAccumUnit/ReadPipeline/RemapCache/RemapCache.sv"
`include "TileAccumUnit/ReadPipeline/Allocator.sv"
`include "TileAccumUnit/ReadPipeline/SramWriteCollector.sv"
`include "TileAccumUnit/ReadPipeline/ReadPipeline.sv"
