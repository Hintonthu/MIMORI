`include "define.sv"
`include "common/SRAM.sv"
`include "common/Semaphore.sv"
`include "common/ND.sv"
`include "common/BitOperation.sv"
`include "common/Controllers.sv"
`include "common/Registers.sv"
`include "common/OffsetStage.sv"
`include "TileAccumUnit/common/OrCrossBar.sv"
`include "TileAccumUnit/common/BofsExpand.sv"
`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooperIndexStage.sv"
`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooperStencilStage.sv"
`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooperMemofsStage.sv"
`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooperVectorStage.sv"
`include "TileAccumUnit/common/AccumWarpLooper.sv"
`include "TileAccumUnit/AccumBlockLooper.sv"
`include "TileAccumUnit/AluPipeline/Simd/Alu.sv"
`include "TileAccumUnit/AluPipeline/Simd/SimdDriver.sv"
`include "TileAccumUnit/AluPipeline/Simd/SimdOperand.sv"
`include "TileAccumUnit/AluPipeline/Simd/SimdTmpBuffer.sv"
`include "TileAccumUnit/AluPipeline/Simd.sv"
`include "TileAccumUnit/AluPipeline/AluPipeline.sv"
`include "TileAccumUnit/WritePipeline/DramWriteCollector/DramWriteCollectorAddrDecode.sv"
`include "TileAccumUnit/WritePipeline/DramWriteCollector/DramWriteCollectorOutput.sv"
`include "TileAccumUnit/WritePipeline/DramWriteCollector.sv"
`include "TileAccumUnit/WritePipeline/WritePipeline.sv"
`include "TileAccumUnit/ReadPipeline/RemapCache/BankSramReadIf.sv"
`include "TileAccumUnit/ReadPipeline/RemapCache/BankSramWriteButterflyIf.sv"
`include "TileAccumUnit/ReadPipeline/RemapCache/RemapCache.sv"
`include "TileAccumUnit/ReadPipeline/Allocator.sv"
`include "TileAccumUnit/ReadPipeline/ChunkAddrLooper/ChunkRowStart.sv"
`include "TileAccumUnit/ReadPipeline/ChunkAddrLooper/ChunkRow.sv"
`include "TileAccumUnit/ReadPipeline/ChunkAddrLooper.sv"
`include "TileAccumUnit/ReadPipeline/ChunkHead.sv"
`include "TileAccumUnit/ReadPipeline/LinearCollector.sv"
`include "TileAccumUnit/ReadPipeline/SramWriteCollector.sv"
`include "TileAccumUnit/ReadPipeline/ReadPipeline.sv"
`include "TileAccumUnit/DramArbiter.sv"
`include "TileAccumUnit/TileAccumUnit.sv"
`include "ParallelBlockLooper.sv"
`include "Top.sv"
