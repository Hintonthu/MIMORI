`include "define.sv"
`include "common/ND.sv"
`include "common/BitOperation.sv"
`include "common/Controllers.sv"
`include "common/Registers.sv"
`include "common/OffsetStage.sv"
`include "common/IndexStage.sv"
`include "common/MemofsStage.sv"
`include "TileAccumUnit/common/AccumBlockLooper.sv"
