`include "define.sv"
`include "common/SRAM.sv"
`include "common/ND.sv"
`include "common/BitOperation.sv"
`include "common/Controllers.sv"
`include "common/OffsetStage.sv"
`include "common/Semaphore.sv"
`include "TileAccumUnit/common/BofsExpand.sv"
`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooperIndexStage.sv"
`include "TileAccumUnit/AluPipeline/Simd/Alu.sv"
`include "TileAccumUnit/AluPipeline/Simd/SimdDriver.sv"
`include "TileAccumUnit/AluPipeline/Simd/SimdOperand.sv"
`include "TileAccumUnit/AluPipeline/Simd/SimdTmpBuffer.sv"
`include "TileAccumUnit/AluPipeline/Simd.sv"
`include "TileAccumUnit/AluPipeline/AluPipeline.sv"
