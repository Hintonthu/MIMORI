`include "TileAccumUnit/WritePipeline/DramWriteCollector/DramWriteCollector.sv"
