`include "ParallelBlockLooper_mc.sv"
