`include "TileAccumUnit/AluPipeline/AluPipeline.sv"
