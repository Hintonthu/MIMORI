`include "TileAccumUnit/ReadPipeline/ReadPipeline_sd.sv"
