`include "TileAccumUnit/ReadPipeline/Allocator.sv"
