`include "define.sv"
`include "common/ND.sv"
`include "common/BitOperation.sv"
`include "common/Controllers.sv"
`include "common/Registers.sv"
`include "common/OffsetStage.sv"
`include "common/IndexStage.sv"
`include "common/MemofsStage.sv"
`include "TileAccumUnit/common/OrCrossBar.sv"
`include "TileAccumUnit/common/AccumBlockLooper.sv"
`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooperCollector.sv"
`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooperIndexStage.sv"
`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooperMemofsStage.sv"
`include "TileAccumUnit/common/AccumWarpLooper/AccumWarpLooperVectorStage.sv"
`include "TileAccumUnit/common/AccumWarpLooper.sv"
`include "TileAccumUnit/WritePipeline/DramWriteCollector/DramWriteCollectorAddrDecode.sv"
`include "TileAccumUnit/WritePipeline/DramWriteCollector/DramWriteCollectorOutput.sv"
`include "TileAccumUnit/WritePipeline/DramWriteCollector.sv"
`include "TileAccumUnit/WritePipeline/WritePipeline.sv"
