`include "TileAccumUnit/DmaPipeline/ChunkAddrLooper/ChunkAddrLooper.sv"
