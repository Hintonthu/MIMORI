`include "Top.sv"
